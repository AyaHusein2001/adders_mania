/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Mon Oct 31 18:23:41 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3864487568 */

module full_adder__0_40(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(o_sum));
endmodule

module full_adder__0_44(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_48(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_52(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_56(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_60(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_64(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_68(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_72(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_76(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_80(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_84(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_88(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_92(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_96(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_100(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_104(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_108(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_112(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_116(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_120(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_124(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_128(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_132(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_136(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_140(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_144(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_148(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_152(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_156(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_160(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module carry_lookahead_adder_32_bit(i_add1, i_add2, o_result, cout, OF);
   input [31:0]i_add1;
   input [31:0]i_add2;
   output [31:0]o_result;
   output cout;
   output OF;

   wire n_0_0_0;
   wire n_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_1;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_2;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_3;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_4;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_5;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_6;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_7;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_8;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_9;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_10;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_11;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_12;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_13;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_14;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_15;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_16;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_17;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_18;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_19;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_20;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_21;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_22;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_23;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_24;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_25;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_26;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_27;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_28;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_29;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire w_G;
   wire n_0_0_63;

   full_adder__0_40 genblk1_0_adderlook (.i_bit1(i_add1[0]), .i_bit2(i_add2[0]), 
      .i_carry(), .o_sum(o_result[0]), .o_carry());
   full_adder__0_44 genblk1_1_adderlook (.i_bit1(i_add1[1]), .i_bit2(i_add2[1]), 
      .i_carry(w_G), .o_sum(o_result[1]), .o_carry());
   full_adder__0_48 genblk1_2_adderlook (.i_bit1(i_add1[2]), .i_bit2(i_add2[2]), 
      .i_carry(n_0_29), .o_sum(o_result[2]), .o_carry());
   full_adder__0_52 genblk1_3_adderlook (.i_bit1(i_add1[3]), .i_bit2(i_add2[3]), 
      .i_carry(n_0_28), .o_sum(o_result[3]), .o_carry());
   full_adder__0_56 genblk1_4_adderlook (.i_bit1(i_add1[4]), .i_bit2(i_add2[4]), 
      .i_carry(n_0_27), .o_sum(o_result[4]), .o_carry());
   full_adder__0_60 genblk1_5_adderlook (.i_bit1(i_add1[5]), .i_bit2(i_add2[5]), 
      .i_carry(n_0_26), .o_sum(o_result[5]), .o_carry());
   full_adder__0_64 genblk1_6_adderlook (.i_bit1(i_add1[6]), .i_bit2(i_add2[6]), 
      .i_carry(n_0_25), .o_sum(o_result[6]), .o_carry());
   full_adder__0_68 genblk1_7_adderlook (.i_bit1(i_add1[7]), .i_bit2(i_add2[7]), 
      .i_carry(n_0_24), .o_sum(o_result[7]), .o_carry());
   full_adder__0_72 genblk1_8_adderlook (.i_bit1(i_add1[8]), .i_bit2(i_add2[8]), 
      .i_carry(n_0_23), .o_sum(o_result[8]), .o_carry());
   full_adder__0_76 genblk1_9_adderlook (.i_bit1(i_add1[9]), .i_bit2(i_add2[9]), 
      .i_carry(n_0_22), .o_sum(o_result[9]), .o_carry());
   full_adder__0_80 genblk1_10_adderlook (.i_bit1(i_add1[10]), .i_bit2(
      i_add2[10]), .i_carry(n_0_21), .o_sum(o_result[10]), .o_carry());
   full_adder__0_84 genblk1_11_adderlook (.i_bit1(i_add1[11]), .i_bit2(
      i_add2[11]), .i_carry(n_0_20), .o_sum(o_result[11]), .o_carry());
   full_adder__0_88 genblk1_12_adderlook (.i_bit1(i_add1[12]), .i_bit2(
      i_add2[12]), .i_carry(n_0_19), .o_sum(o_result[12]), .o_carry());
   full_adder__0_92 genblk1_13_adderlook (.i_bit1(i_add1[13]), .i_bit2(
      i_add2[13]), .i_carry(n_0_18), .o_sum(o_result[13]), .o_carry());
   full_adder__0_96 genblk1_14_adderlook (.i_bit1(i_add1[14]), .i_bit2(
      i_add2[14]), .i_carry(n_0_17), .o_sum(o_result[14]), .o_carry());
   full_adder__0_100 genblk1_15_adderlook (.i_bit1(i_add1[15]), .i_bit2(
      i_add2[15]), .i_carry(n_0_16), .o_sum(o_result[15]), .o_carry());
   full_adder__0_104 genblk1_16_adderlook (.i_bit1(i_add1[16]), .i_bit2(
      i_add2[16]), .i_carry(n_0_15), .o_sum(o_result[16]), .o_carry());
   full_adder__0_108 genblk1_17_adderlook (.i_bit1(i_add1[17]), .i_bit2(
      i_add2[17]), .i_carry(n_0_14), .o_sum(o_result[17]), .o_carry());
   full_adder__0_112 genblk1_18_adderlook (.i_bit1(i_add1[18]), .i_bit2(
      i_add2[18]), .i_carry(n_0_13), .o_sum(o_result[18]), .o_carry());
   full_adder__0_116 genblk1_19_adderlook (.i_bit1(i_add1[19]), .i_bit2(
      i_add2[19]), .i_carry(n_0_12), .o_sum(o_result[19]), .o_carry());
   full_adder__0_120 genblk1_20_adderlook (.i_bit1(i_add1[20]), .i_bit2(
      i_add2[20]), .i_carry(n_0_11), .o_sum(o_result[20]), .o_carry());
   full_adder__0_124 genblk1_21_adderlook (.i_bit1(i_add1[21]), .i_bit2(
      i_add2[21]), .i_carry(n_0_10), .o_sum(o_result[21]), .o_carry());
   full_adder__0_128 genblk1_22_adderlook (.i_bit1(i_add1[22]), .i_bit2(
      i_add2[22]), .i_carry(n_0_9), .o_sum(o_result[22]), .o_carry());
   full_adder__0_132 genblk1_23_adderlook (.i_bit1(i_add1[23]), .i_bit2(
      i_add2[23]), .i_carry(n_0_8), .o_sum(o_result[23]), .o_carry());
   full_adder__0_136 genblk1_24_adderlook (.i_bit1(i_add1[24]), .i_bit2(
      i_add2[24]), .i_carry(n_0_7), .o_sum(o_result[24]), .o_carry());
   full_adder__0_140 genblk1_25_adderlook (.i_bit1(i_add1[25]), .i_bit2(
      i_add2[25]), .i_carry(n_0_6), .o_sum(o_result[25]), .o_carry());
   full_adder__0_144 genblk1_26_adderlook (.i_bit1(i_add1[26]), .i_bit2(
      i_add2[26]), .i_carry(n_0_5), .o_sum(o_result[26]), .o_carry());
   full_adder__0_148 genblk1_27_adderlook (.i_bit1(i_add1[27]), .i_bit2(
      i_add2[27]), .i_carry(n_0_4), .o_sum(o_result[27]), .o_carry());
   full_adder__0_152 genblk1_28_adderlook (.i_bit1(i_add1[28]), .i_bit2(
      i_add2[28]), .i_carry(n_0_3), .o_sum(o_result[28]), .o_carry());
   full_adder__0_156 genblk1_29_adderlook (.i_bit1(i_add1[29]), .i_bit2(
      i_add2[29]), .i_carry(n_0_2), .o_sum(o_result[29]), .o_carry());
   full_adder__0_160 genblk1_30_adderlook (.i_bit1(i_add1[30]), .i_bit2(
      i_add2[30]), .i_carry(n_0_1), .o_sum(o_result[30]), .o_carry());
   full_adder genblk1_31_adderlook (.i_bit1(i_add1[31]), .i_bit2(i_add2[31]), 
      .i_carry(n_0_0), .o_sum(o_result[31]), .o_carry());
   NAND2_X1 i_0_0_0 (.A1(n_0_0_62), .A2(n_0_0_0), .ZN(cout));
   OAI21_X1 i_0_0_1 (.A(n_0_0), .B1(i_add1[31]), .B2(i_add2[31]), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_2 (.A1(n_0_0_2), .A2(n_0_0_1), .ZN(n_0_0));
   OAI21_X1 i_0_0_3 (.A(n_0_1), .B1(i_add1[30]), .B2(i_add2[30]), .ZN(n_0_0_1));
   NAND2_X1 i_0_0_4 (.A1(i_add2[30]), .A2(i_add1[30]), .ZN(n_0_0_2));
   NAND2_X1 i_0_0_5 (.A1(n_0_0_4), .A2(n_0_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_0_6 (.A1(i_add2[29]), .A2(i_add1[29]), .ZN(n_0_0_3));
   OAI21_X1 i_0_0_7 (.A(n_0_2), .B1(i_add1[29]), .B2(i_add2[29]), .ZN(n_0_0_4));
   NAND2_X1 i_0_0_8 (.A1(n_0_0_6), .A2(n_0_0_5), .ZN(n_0_2));
   OAI21_X1 i_0_0_9 (.A(n_0_3), .B1(i_add1[28]), .B2(i_add2[28]), .ZN(n_0_0_5));
   NAND2_X1 i_0_0_10 (.A1(i_add2[28]), .A2(i_add1[28]), .ZN(n_0_0_6));
   NAND2_X1 i_0_0_11 (.A1(n_0_0_8), .A2(n_0_0_7), .ZN(n_0_3));
   NAND2_X1 i_0_0_12 (.A1(i_add2[27]), .A2(i_add1[27]), .ZN(n_0_0_7));
   OAI21_X1 i_0_0_13 (.A(n_0_4), .B1(i_add1[27]), .B2(i_add2[27]), .ZN(n_0_0_8));
   NAND2_X1 i_0_0_14 (.A1(n_0_0_10), .A2(n_0_0_9), .ZN(n_0_4));
   OAI21_X1 i_0_0_15 (.A(n_0_5), .B1(i_add1[26]), .B2(i_add2[26]), .ZN(n_0_0_9));
   NAND2_X1 i_0_0_16 (.A1(i_add2[26]), .A2(i_add1[26]), .ZN(n_0_0_10));
   NAND2_X1 i_0_0_17 (.A1(n_0_0_12), .A2(n_0_0_11), .ZN(n_0_5));
   NAND2_X1 i_0_0_18 (.A1(i_add2[25]), .A2(i_add1[25]), .ZN(n_0_0_11));
   OAI21_X1 i_0_0_19 (.A(n_0_6), .B1(i_add1[25]), .B2(i_add2[25]), .ZN(n_0_0_12));
   NAND2_X1 i_0_0_20 (.A1(n_0_0_14), .A2(n_0_0_13), .ZN(n_0_6));
   OAI21_X1 i_0_0_21 (.A(n_0_7), .B1(i_add1[24]), .B2(i_add2[24]), .ZN(n_0_0_13));
   NAND2_X1 i_0_0_22 (.A1(i_add2[24]), .A2(i_add1[24]), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_23 (.A1(n_0_0_16), .A2(n_0_0_15), .ZN(n_0_7));
   NAND2_X1 i_0_0_24 (.A1(i_add2[23]), .A2(i_add1[23]), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_25 (.A(n_0_8), .B1(i_add1[23]), .B2(i_add2[23]), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_26 (.A1(n_0_0_18), .A2(n_0_0_17), .ZN(n_0_8));
   OAI21_X1 i_0_0_27 (.A(n_0_9), .B1(i_add1[22]), .B2(i_add2[22]), .ZN(n_0_0_17));
   NAND2_X1 i_0_0_28 (.A1(i_add2[22]), .A2(i_add1[22]), .ZN(n_0_0_18));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_20), .A2(n_0_0_19), .ZN(n_0_9));
   NAND2_X1 i_0_0_30 (.A1(i_add2[21]), .A2(i_add1[21]), .ZN(n_0_0_19));
   OAI21_X1 i_0_0_31 (.A(n_0_10), .B1(i_add1[21]), .B2(i_add2[21]), .ZN(n_0_0_20));
   NAND2_X1 i_0_0_32 (.A1(n_0_0_22), .A2(n_0_0_21), .ZN(n_0_10));
   OAI21_X1 i_0_0_33 (.A(n_0_11), .B1(i_add1[20]), .B2(i_add2[20]), .ZN(n_0_0_21));
   NAND2_X1 i_0_0_34 (.A1(i_add2[20]), .A2(i_add1[20]), .ZN(n_0_0_22));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_24), .A2(n_0_0_23), .ZN(n_0_11));
   NAND2_X1 i_0_0_36 (.A1(i_add2[19]), .A2(i_add1[19]), .ZN(n_0_0_23));
   OAI21_X1 i_0_0_37 (.A(n_0_12), .B1(i_add1[19]), .B2(i_add2[19]), .ZN(n_0_0_24));
   NAND2_X1 i_0_0_38 (.A1(n_0_0_26), .A2(n_0_0_25), .ZN(n_0_12));
   OAI21_X1 i_0_0_39 (.A(n_0_13), .B1(i_add1[18]), .B2(i_add2[18]), .ZN(n_0_0_25));
   NAND2_X1 i_0_0_40 (.A1(i_add2[18]), .A2(i_add1[18]), .ZN(n_0_0_26));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_28), .A2(n_0_0_27), .ZN(n_0_13));
   NAND2_X1 i_0_0_42 (.A1(i_add2[17]), .A2(i_add1[17]), .ZN(n_0_0_27));
   OAI21_X1 i_0_0_43 (.A(n_0_14), .B1(i_add1[17]), .B2(i_add2[17]), .ZN(n_0_0_28));
   NAND2_X1 i_0_0_44 (.A1(n_0_0_30), .A2(n_0_0_29), .ZN(n_0_14));
   OAI21_X1 i_0_0_45 (.A(n_0_15), .B1(i_add1[16]), .B2(i_add2[16]), .ZN(n_0_0_29));
   NAND2_X1 i_0_0_46 (.A1(i_add2[16]), .A2(i_add1[16]), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_47 (.A1(n_0_0_32), .A2(n_0_0_31), .ZN(n_0_15));
   NAND2_X1 i_0_0_48 (.A1(i_add2[15]), .A2(i_add1[15]), .ZN(n_0_0_31));
   OAI21_X1 i_0_0_49 (.A(n_0_16), .B1(i_add1[15]), .B2(i_add2[15]), .ZN(n_0_0_32));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_34), .A2(n_0_0_33), .ZN(n_0_16));
   OAI21_X1 i_0_0_51 (.A(n_0_17), .B1(i_add1[14]), .B2(i_add2[14]), .ZN(n_0_0_33));
   NAND2_X1 i_0_0_52 (.A1(i_add2[14]), .A2(i_add1[14]), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_53 (.A1(n_0_0_36), .A2(n_0_0_35), .ZN(n_0_17));
   NAND2_X1 i_0_0_54 (.A1(i_add2[13]), .A2(i_add1[13]), .ZN(n_0_0_35));
   OAI21_X1 i_0_0_55 (.A(n_0_18), .B1(i_add1[13]), .B2(i_add2[13]), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_56 (.A1(n_0_0_38), .A2(n_0_0_37), .ZN(n_0_18));
   OAI21_X1 i_0_0_57 (.A(n_0_19), .B1(i_add1[12]), .B2(i_add2[12]), .ZN(n_0_0_37));
   NAND2_X1 i_0_0_58 (.A1(i_add2[12]), .A2(i_add1[12]), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_40), .A2(n_0_0_39), .ZN(n_0_19));
   NAND2_X1 i_0_0_60 (.A1(i_add2[11]), .A2(i_add1[11]), .ZN(n_0_0_39));
   OAI21_X1 i_0_0_61 (.A(n_0_20), .B1(i_add1[11]), .B2(i_add2[11]), .ZN(n_0_0_40));
   NAND2_X1 i_0_0_62 (.A1(n_0_0_42), .A2(n_0_0_41), .ZN(n_0_20));
   OAI21_X1 i_0_0_63 (.A(n_0_21), .B1(i_add1[10]), .B2(i_add2[10]), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_64 (.A1(i_add2[10]), .A2(i_add1[10]), .ZN(n_0_0_42));
   NAND2_X1 i_0_0_65 (.A1(n_0_0_44), .A2(n_0_0_43), .ZN(n_0_21));
   NAND2_X1 i_0_0_66 (.A1(i_add2[9]), .A2(i_add1[9]), .ZN(n_0_0_43));
   OAI21_X1 i_0_0_67 (.A(n_0_22), .B1(i_add1[9]), .B2(i_add2[9]), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_46), .A2(n_0_0_45), .ZN(n_0_22));
   OAI21_X1 i_0_0_69 (.A(n_0_23), .B1(i_add1[8]), .B2(i_add2[8]), .ZN(n_0_0_45));
   NAND2_X1 i_0_0_70 (.A1(i_add2[8]), .A2(i_add1[8]), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_48), .A2(n_0_0_47), .ZN(n_0_23));
   NAND2_X1 i_0_0_72 (.A1(i_add2[7]), .A2(i_add1[7]), .ZN(n_0_0_47));
   OAI21_X1 i_0_0_73 (.A(n_0_24), .B1(i_add1[7]), .B2(i_add2[7]), .ZN(n_0_0_48));
   NAND2_X1 i_0_0_74 (.A1(n_0_0_50), .A2(n_0_0_49), .ZN(n_0_24));
   OAI21_X1 i_0_0_75 (.A(n_0_25), .B1(i_add1[6]), .B2(i_add2[6]), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_76 (.A1(i_add2[6]), .A2(i_add1[6]), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_77 (.A1(n_0_0_52), .A2(n_0_0_51), .ZN(n_0_25));
   NAND2_X1 i_0_0_78 (.A1(i_add2[5]), .A2(i_add1[5]), .ZN(n_0_0_51));
   OAI21_X1 i_0_0_79 (.A(n_0_26), .B1(i_add1[5]), .B2(i_add2[5]), .ZN(n_0_0_52));
   NAND2_X1 i_0_0_80 (.A1(n_0_0_54), .A2(n_0_0_53), .ZN(n_0_26));
   OAI21_X1 i_0_0_81 (.A(n_0_27), .B1(i_add1[4]), .B2(i_add2[4]), .ZN(n_0_0_53));
   NAND2_X1 i_0_0_82 (.A1(i_add2[4]), .A2(i_add1[4]), .ZN(n_0_0_54));
   NAND2_X1 i_0_0_83 (.A1(n_0_0_56), .A2(n_0_0_55), .ZN(n_0_27));
   NAND2_X1 i_0_0_84 (.A1(i_add2[3]), .A2(i_add1[3]), .ZN(n_0_0_55));
   OAI21_X1 i_0_0_85 (.A(n_0_28), .B1(i_add1[3]), .B2(i_add2[3]), .ZN(n_0_0_56));
   NAND2_X1 i_0_0_86 (.A1(n_0_0_58), .A2(n_0_0_57), .ZN(n_0_28));
   OAI21_X1 i_0_0_87 (.A(n_0_29), .B1(i_add1[2]), .B2(i_add2[2]), .ZN(n_0_0_57));
   NAND2_X1 i_0_0_88 (.A1(i_add2[2]), .A2(i_add1[2]), .ZN(n_0_0_58));
   NOR2_X1 i_0_0_89 (.A1(n_0_0_60), .A2(n_0_0_59), .ZN(n_0_29));
   NOR2_X1 i_0_0_90 (.A1(i_add1[1]), .A2(w_G), .ZN(n_0_0_59));
   AOI21_X1 i_0_0_91 (.A(i_add2[1]), .B1(i_add1[1]), .B2(w_G), .ZN(n_0_0_60));
   OAI22_X1 i_0_0_92 (.A1(n_0_0_61), .A2(i_add2[31]), .B1(n_0_0_62), .B2(
      o_result[31]), .ZN(OF));
   NAND2_X1 i_0_0_93 (.A1(n_0_0_63), .A2(o_result[31]), .ZN(n_0_0_61));
   NAND2_X1 i_0_0_94 (.A1(i_add2[31]), .A2(i_add1[31]), .ZN(n_0_0_62));
   AND2_X1 i_0_0_95 (.A1(i_add2[0]), .A2(i_add1[0]), .ZN(w_G));
   INV_X1 i_0_0_96 (.A(i_add1[31]), .ZN(n_0_0_63));
endmodule
